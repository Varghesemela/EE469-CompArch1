module Decoder(input [4:0] write_reg, 
               input Regwrite, 
               output write_en)
